// See LICENSE for license details.
module AdderExtModule(
  input [15:0] foo,
  output [15:0] bar
);
  assign bar = foo + 1;
endmodule

