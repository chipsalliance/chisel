module BlackBoxPassthrough2(
    input  [0:0] in,
    output [0:0] out
);
  assign out = in;
endmodule
