
module SimpleExtModule(
  input [15:0] foo,
  output [15:0] bar
);
  assign bar = foo;
endmodule

