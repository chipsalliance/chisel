module ExtPath(); endmodule
