// SPDX-License-Identifier: Apache-2.0
`ifndef _parameters_vh_
`define _parameters_vh_
parameter VALUE = 2;
`endif
