// See LICENSE for license details.
`ifndef _parameters_vh_
`define _parameters_vh_
parameter VALUE = 2;
`endif
